-- https://allaboutfpga.com/vhdl-4-to-1-mux-multiplexer/
--https://steemit.com/logic/@drifter1/logic-design-vhdl-basic-circuits


library IEEE;
use IEEE.std_logic_164.all;

entity mux_4to1 is
    port(
        A, B, C, D  :   in std_logic;
        S0, S1          :   in std_logic;
        Z               :   out std_logic
    );
end mux_4to1;

architecture behavior of mux_4to1 is
begin
process (A, B, C, D, S0, S1) is
    begin
        Z <= A when S1='0' and S0='0' else
             B when S1='0' and S0='1' else
             C when S1='1' and S0='0' else
            when S1='1' and S0='1';
end process;
end behavior;


-- testbench for mux
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY tb_mux IS
END tb_mux;
 
ARCHITECTURE behavior OF tb_mux IS
 
    – Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT mux_4to1
    PORT(
         A : IN  std_logic;
         B : IN  std_logic;
         C : IN  std_logic;
         D : IN  std_logic;
         S0 : IN  std_logic;
         S1 : IN  std_logic;
         Z : OUT  std_logic
        );
    END COMPONENT;
 
   – Inputs
   signal A : std_logic := '0';
   signal B : std_logic := '0';
   signal C : std_logic := '0';
   signal D : std_logic := '0';
   signal S0 : std_logic := '0';
   signal S1 : std_logic := '0';
 
    --Outputs
   signal Z : std_logic;
 
BEGIN
 
     – Instantiate the Unit Under Test (UUT)
   uut: mux_4to1 PORT MAP (
          A => A,
          B => B,
          C => C,
          D => D,
          S0 => S0,
          S1 => S1,
          Z => Z
        );
 
   – Stimulus process
   stim_proc: process
   begin
      – hold reset state for 100 ns.
      wait for 100 ns; 
 
    A <= '1';
    B <= '0';
    C <= '1';
    D <= '0';       
 
    S0 <= '0'; S1 <= '0';
 
      wait for 100 ns; 
 
    S0 <= '1'; S1 <= '0';
 
      wait for 100 ns; 
 
    S0 <= '0'; S1 <= '1';
 
        wait for 100 ns;   
 
    S0 <= '0'; S1 <= '1';  
 
        wait for 100 ns;   
 
    end process;
 
END;
